class f_sequence_item extends uvm_sequence_item;
  rand bit i_wren;
  rand bit i_rden;
  rand bit [7:0] i_wdata;
  bit full;
  bit empty;
  bit o_alm_full;
  bit o_alm_empty;
  bit [7:0] o_rdata;
  
  `uvm_object_utils_begin(f_sequence_item)
  `uvm_field_int(i_wren, UVM_ALL_ON)
  `uvm_field_int(i_rden, UVM_ALL_ON)
  `uvm_field_int(i_wdata, UVM_ALL_ON)
  `uvm_object_utils_end
  constraint wr_rd2 {wr != rd;}
  
  function new(string name = "f_sequence_item");
    super.new(name);
  endfunction

endclass
